// This is the EX/MEM pipeline register
module EX_MEM_reg
(
    clk,
    rst,
);

    input clk, rst;

endmodule
