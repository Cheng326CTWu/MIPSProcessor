// This is the ID/EX pipeline register
module ID_EX_reg
(
    clk,
    rst,
);

    input clk, rst;

endmodule
