// This is the MEM/WB pipeline register
module MEM_WB_reg
(
    clk,
    rst,
);

    input clk, rst;

endmodule
